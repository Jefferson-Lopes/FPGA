��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��L�+�h�0I��y�������b�~�L�ʬ3�&�;��eW����x�k�Ր�7\�?^ �R����:�{|�h.9��4!�B~����/!���o_mnKD��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:��WJ}KV��g���ơH-��I�g�E�w�/)
�_�{Ei)��p6���Ϳ��µ���I��j���*�:��f�)��yP�d�VAm�
Tȧ��S�cfrY�b'�.����Z�Q��[R���h�Ȧ�d��Q���V�� 9��$����'A��ũ�i�'�ߵ��1����-T%~T�)A`�2�����B�DM�9�'��f[�P�zj]�4���R�mN��)8��MÇ�()٬�=�����u�(� x>\A�
\p�ԁ�5f��궾��l5ş*PZ/1	_nn�U,ɓA���ӛ{�:1<���'��~y�����sA����WJ��q5��-���ԅ�Y���Rta�ǒ�M.���{�������-@:?�O�z�f~84R5J������dí����D�БP�@���ҩc'�JՏ�Q�H���}��W�`ƵX��*�`&Q����(;ǴBZ���zo����(����=%��=Ed�$�޸;ku�[|�25��o�BOrA?8�����b���1�`K�T�,�P��c�.`h:�|��"�Ӆ�b�?�� c�,(h��_��#�$$���ED���:K����m/i���j���Uh54,a!����^��w>)ׂ�ϭ��^�/3L�8:���$6���%�*sl�����~'�p�&�R�Q�;d�T�p��\7�m�S|v�ql��'%�S��v��I�N�j�A��$;`6��j-ac�LW��O<�|���ЂhUD'���4C�Vu�[X$��H"R>X��5�4=�����ÙOQ��z<�f�Zjq�/��.<rx�-GX(@`~$r%Ԯ�Es�9��h.f�S���7__��Y���r�K�L#v�����+n� =�
!�G�>�[x�����xD1��D�'|�q����d�`�Wjk��X�1US��Ѭ(i
HB�v�{eͅ��z.%���O����E>2�������a�Dľv�B����"�����;t�����3��HF�ԛ8	]*��x���Xz��xZ�]*��"( ���z�ecn��)>M��Z2�_+��@(���6Y��M��
���\��ĉ�Dǲ�O�h�f�Y� �~��Z��1ܜ�� �9�_S����y��Y��E����<���g;-�Ew��Ve�},"��)�(6\����j'��&]K������Wx.�z��Ο����i�Ulh���J�0+6������m������\7�ܘ(N��p��P�����Y`�o���+`D�8��q��#���5hO5�)}���@�le���^�]�k�Y}	D�H"*�����})����I3��E3�K'��g<jc��Ƿgr�K$��>�q�����Ξ E�[�w��K��mb��?���v��*ƿ��8���� #��4�.Zl�l1k4���e��@H�5��múF��#�� �kY�o���d���Ga��.��L��|�CG�C�*tp�X�)7�技�K!eŮ���H4j��	h�M�.�|Bk��K�C�q�Z�ߤK���X�/O�[���@��QW+t����}��..�����4`��D���_�5�*�i���UԔ��&���� 8���G��-����zc��H˔̅H�!>-ݏ�ݩ��F���}]���A��Vr��������	����Q/��/���n��+\J&�,��7�����N��j��Z� eR9'��dK�s/���$�Ԗ��!��Z��!z��?��ǅ�F�W�h����;�9׷���Q�>P%�*$��	���x@�$�K�W#$���G�qP�ݟҹ �1��|������*�G����F�e ��]=$g&��%,x,�>z��G{X�FA)B&h�u���^�Y�5���vC���� ��Y�:K%���-�(�kR��f�"��r5��&��
��/\�l^D�ɹ�9����]��i�L���xoU�W^uyD\�3[	�~�d�)�:�O#��F���Oy��o4�|���fU�t=4��J����o���Wt6� �]���W1�w���x� ��;�-�׫ʫ�.���PZƊO�F���
��^n}t�Xuud��e�B��������D`B����ΩeZ��d��[�����
�z<(	-񋮰�!�Xi�g����l�� ����	��&�`3��B8���P���P��M�*ZS^�v_|���kJQr�k��Z��3_��#	�im!?��}K�i� '�Qm13~�z,�Z3�B�h���S�7�$�]�k�DV��9d G�����@�1����z� 7�x YL�X��l�X�W�p_��Ppik���W�oH�tB��Ӳ��ms!-��.��s�74�·�Zɕ(gz�.f��ǁA���P����:Lv7��DA�9�X��1��MY���|�6'��8��B( ��"���	�� 9�f�?
T��C��γ]�B�U�8�3�i���1�Q$���D&�4$�����!�h˾[��.����TN�>��;��ʈ�"<Ʋ/�k��A@�r�7ios��\�|F�>�;���0=����1��jJ;�.�p����~��_�����Rre
w^��'��O-GoV窍fX����}ߦ8'�����έ�ZfG�����QA���>�_�!*�6���4sϦ�J[�
DX�_�Cs��<��V��($b��9�+�՟9�>h���A�.���[Y9�	����."Q"���A-TH�i��q��2*�k������e���f4@���() ���0��k�x��܀ Ӕ�7 V�0�;T�m ���<C�o�2�)�ej2����ל�m)��������7e����9�mі2������2m�.I�9������S�u�0�}��L��_�	a�C��}��|�a����@֗3��3��L0`/ܜ��v�����tr'm�ƕ�����ר?n'�k�ݜ�GjAL���8� ����n��5��b������:�Zh���ȥ��ܹ���a&�Fw��\P�\��B�aIC�0�q��ѹ�@����+�|b�9�-���R�:���T�R&LH[��b����ӯ��@@Z� `���u8��^�e���)�綉ZZ3��/��P}>�x�9�0�{����l�݋xk��������l��c�̴U���N\p@�~�.á����OOv�<f�u�ӵY���F�+pVɝ&L�tՃ�]����Q����"��ƽ�b3fEVa��UoTW�%�#�AQ�>8�e�b@�'�l)���7��l�L��}_B�\
dG�i���L�g�,��Ү*�����[��Q|�������u�s�R�`E9BPǘi��?.ֳ*���a����@�~T��ӵ^+>�"S#u�6�+��2��Y������[tH(���Y}�%�ߜ4	��H"E�?���c63���f�s���Խ=�ǆ.Ci�u�'�Ӆj�]�������{��x6H*�  ���{���BxZ��B)��ñ�[�A5��8k_�Է���}��`�����Ȟ.U�>V���M��;psKSQ�	���d�lO(z���4���Κ?zKx=:ԗ�q�B}sU��v���=��v���6�Π?��P+,bYr�8������gL�nS�٨��)�U�ll5Ȟ�q���R��,D�Dv��V�"-�+o�P$������4O��I�aOTa�i��Yc'5鋂�)�*����P$�dy�-[�,)۩�¬[�F�R�ó#�w&&l�ty̅M����*��j%$�\A��ngp�?����V+�b~�oB��ʧsv�Qz�P	�SlS#9F�O"K�k霍���]��q�遺ib]��o�`�~�}^/#_Sp]c��⦍���7V�Ʊ���	v��}����a(1�䴃�>`dk�i''�9��ܠ�6
�U�o���D�[�`���5�]��Vz��{=J���2C%��6��Ż�t�B#��w�)3��⁤���:��� �@���Nc�Q:p��%�Wx��O���I8�T|!��wg�܌�M�s������$�,��Ron�#��Y�Ò%���������H��=8ioO5P
���؉��&���[�*�@�����?��,o�:�f&�䐋7v}	@�����y�m�.���z^tQ~Ow$=��"�摩j$,}7�L��>�c�n�c����6����8P�q�%�X"��&9	p�}#Q��Q���M���(}�d����A�iۆ������̵�"L �(�ȥ�>�SH���I�]�Cb��YHW:�P2���I;%�l c>y��V���h(�2��AUX#�l�C�� y��� �y�)0�9M��p�5��aR�~[b�0hz��a��r��89���Ex?;�^�ѻ��}�����*j{*�O� kOd1�t�Z^�����-�W�~�Q�[��l��*W�h��K��}[P��}���+YH�S%����Py�8%B��l*����:{�u�X��y�z4�J�l�����\�7�����N��V j�wIg�sgXe*���.E�_/�D��Y���@�UqR���8�H5��q�!�nϻ�X�A��]g�tF����[|��?Px'ҝ���|�SD^<��s�V��~}�ъ����q�C���7k��U��n�򴓊a�!:P����t��;��-�)�*�t��뚴u �� Q�����ˋ�����0U˨=��')���.Ē�,BV���D��[f�}�B�jzi�m�}�5�\N�%-䒰E��� d^�$!�ZuF����O^S�L�Ac\r���Ng/�fe����^I>HUWV\}~D<�.z��4��,������r��z4��I�ו�L�ZM�Xw5$�+�dY+Jw4{eO���g���k��Q����QyKkG?�] X��{�k�Zȃ�윅�E$=�%�����?��}��-��z?$ۚw%}��3���>�!b˦�:��Z#��I����?X�[;\C^��$�殠DCߓ0�T���(�F��,��_�nM, �v ����i�{�a-0"���$"����2@E����dc����rK,d�_�a��%�N��i�!�]�S��� ��ߑ�����'$-.Z��Y����hD�a�	�)�e:ow(���K�5>B�EW"^��ϡ�i}���-4��d�y�� �V��,�z�:�[�[�\���Kb=�o!�њ�ɛRk��ԯT��T�H�4b��]���չO)��h�˪4w�MY�Lx8o�&q���<��Y��^�Lq�;�- ����%��V\���6�D��?�d ���2�
�^�g��J�������˽��H�E� 
/�3x+�R�{/�.*�G��+���7I��2��Uf����&+�՟�E'�|9�Mť�0[ �ӰȀ�(5[U�r��}%!۶��4ލRs@����[�B<�+v�!p�Օ���9N��~ڤ�4�X�i��և�H �M�X'��n��O�� �_^Љ������~�[�ess�J�=x�<���j�J�K0b��9e�d����h�M��Ɲ�y�y
����K����y#�u^���Q��Z�NX(Č�T�-�� E���. �Ği3M�YwAР���� ��z7���u��!����M��$��o����B0fOA�6���ҵj�lX�����S�(���PI�Jp*_V�c��˦�����*\��Z/��3yq|z�gKk���5C�����A��jhm�����_�D��p�Y02����?��!�C�p���A�jX]�}�ڀ]'
��S�"���1����}��%z��@B|�ɸ�wK7�`���倠Tf�����4r�]�z��?]i���Q��\�������E6 e�5N�[�z�n���Kl"lf�+Y÷=(�.X���|�'��s�)��@�SS��F�}��������JGi����&��A � ���5+-��c�dW��������#����Jcp�v*�Ȁ�Zn�N�C�i��3�ܨ��ur�T��	T�����D���^
���g�QA��W�F�{�0�g#���Q<w��[C�'͙W���o`g���sa�D*7�E��iKH������2���3S8�_�!���:�Z���)k��	���Q�?3�3���IRs��
yI2�1ٯ1�zg��K�x�kA����9�@����`�%	�C�WƸ��~#ev���1J\��TB(���������$�D�)���xU��;h�V�i���⿷k�sQ4����A�?hq�r�{|Ru�@ɐY���ܮ�ԇ�ݙNC3DgciC��e��I�e���X��!�d�\K�&�Ϥ��]q�=��#F� ) l�/m�c�[�+1�-�|����ڳ�7��������P��k��.U@䕅���<
^$�L<�!�.�N��ps�e�G�ay�WY�nX�@��|�b��Ys1�'�B�1��':�U��)9��솈�[�>�s�����~x7�ΏMz��Z�`�u�U?m"�pU�;�aj1<���eD�0���qM^*�k���U� y�t�Cǉ"e�@������ⓑ���6Q��"�)0�  *;/8�!:â���yR}>_�U�[6�F��3k�@���㯫�&ci����Z�sp�����[���
e��/�Fٛ���Pr��ѝ��)O�BTF�c��6S�������*��g�>[gy�e�����n�!�ǃ+�Ŝ�|�\B �!�h�ǓP�Kjí�E=Vo��srB��)�g�цYM�d��*}�E�#�.�+�����t��u��7�H��#x8�Ylź���<�O�P,����
}뮣I�æ�i�y��yꡭ�w��J  �a���ݟ�Ͻ�3t�dH��A���?�ғ_+ե�XwӁ�@�%Q���g��V����X��L�YJ�u�Z�Z��1���-APd4�1���Q�9ٿ���*$Y)���Z�4�9pa�������������6E������yd�J�LPa���Vh�'�590�(�N���1;�3ff-1�3�|ʶ�ql=:���1��v�kW2���$�?v2�W��Z(�.NdZ�1Q�۪o�=�ۢ�WQf�/ ����rǘ���|v@�P����iq���,@^uÑ�[&8M���Yl�j*A#�HD��0�����H9G�6ဟ�������*p��A���@Jð�����vݿ�23��e��$�'�p���%Q��X����`�m�*�y]��`�������9ov���sTn5d+��`mz�sЫ$�ĚT�L��X8�
(���r3Ed@��p'�&E�. MĶ�6S�����B�g�֊Al�ҧ��B�xS���T��| ��LDK��$}��ֽPUH�4hЦ5tj���;�����.�ng~7A�>��׫��\�P4���~+���
)���95���9U�G��"�el��L�BFTi_zD��οc*�=bl+|L�q�i���U�1]�k$�9p��8t4�`�#b�:g�F�h]�'�o����,ٛ��$⋯7P����g�M�u�}- ��?�V�!*���0��7���[dl�0�e��G�A��~8.�M��LD���Q 	�*��Ŵ-Z/<�֔��_b�2�(�������}}���U�95�}%42?�=������-s[Ըi���P�`�	��m��R�[��؛P�}��tX̝ߴڑv��N�j4~
�J�N�O�ܭ�9�BM�gg���� ~��IR'^�a�7P~�`�Hi�Dl�/M�$�D�DU6j��M��:��1�N9�� _�A���f�5��oz�G���^+z�� �y�*�MY�A�����Vr�<qNo�9�r�	�xUM)>^�V�+�űn���+y�x�ĩcE������DPm:�x#K0�:�a�%���S�H�n�S��.Sϙz��;�Mt��vK��t{z��)�Ē����N�n�;�>v{��+�4 �]����ՍKٜEsD����,�@ӻQ�l� ��oO��k{,�����J/��R���O�χ��Up�����;>�=)~�=sQ�.`���{P��KU���T���{82��6R�� =|+��Ȩ��f�:�J"�:ʔ8��d����#����`���oZ��кR��������!�+���C�r��p��R8>k���#Z�|8F?l���E�1 ���xp+��S���.J������:���Qއ��d'?͈.k��Tb�]��������=�g��F3���6�6�~ ������dkF2�o$FE/6��@U�g7��a���W�-�Aa����I�~w����
/�w:�Iژ�m>�_E�R|����VȀ�v륒R��bJg�,u�k�	����B�-��������RW�g�߶�*�� 78m������ �<��
�С^z��\}G���Ж��	��9ϐJ����0����_����K4%���7���x����|��(�ǣ|��NN�W[q@�T��@��&~r�	����eNbQ���~�w0��8REǯ��h�HL�~�h�\����P%G��)���eXƾ���jBI�}����:׼�W��g�K��:�ġz�Љ����ڨ�r�5{��
h�n��mB
�ؽlf
4,������Y��4�&UY�O����R�|)��K�l�p��y�qw6O}���u�W,5u�Y����"K�M�����Am������� e�@)���� j��XAk�g�jdpBM�NWYn����3��"6Jn%蛰(E�IÆ��Ǭ|ztdQ��l��D\G0�"�z5)㸛8��F��#��c�8��H�S�_�G�	���&e�Zd��(3&�c��r7�k�(��0^��!������XT��]	s���}~}>��ԣ���d�|��$XY
ǐ�(`��.�f��qQ����{/V·���Ok��L����m��+��7�v%_w[J�����c�,}�0���zoZ��T�X�v�Ix
�j�Vѵ���5b�^y���)wy����ӡ~������K��wЅnе���*	l�]c�Xc���C��'5��&���A2�*c!=�[1�/�۰�g>�>7qh�s��L�͒�;]���$�"� ��z�qr�^�hZe�cd'5�ƀ���I�z<]S�	epW��dn�`E��K>����Z!a�y@ey�Z����ҙ����=_�t�$���f����V�K�^(@j��:S��<�� _{{>ac0��*JSX�ѽg��&�(X�q��$kX��. f������W�أ��w��uC� �J"dWL1/+r��	ܗA�]��S����1q��`��[�X��d'�U�u��Æ��vh�I��h�	���gD���S�R�ߣ�ǣ��� I�\3UtbM�7�s�2t���Is���*,�;���Q�J�Fz��Lok4����y���h�¾m\ST3�wl��F�[q)�V�.�$�睍�����@ӿ(�`�c>�@��_7�9�kNV���6k���2{I��xի�en��u�7���Tf�cS&4�=B�{̽R���u� o�����1P����oz�l"D��Ɍ�4�xr�qè�7"�i�z�O��[\�P���MuP�s��t���ϓ!�Q\b�AJ�!��b3��KQ��@M�>�84��"J��n�#i��'�ATYmѦ�d.���K���WG7�>���S�BzO�q��������f�C?X���K��!�_�P�N|�(�S�K8�V-�t�R�ځ�ݹ�l'�	�,؂]�?-v{�X���0� �� #n)f����
�*a�4���p����^��Wz�]E=0�|��K(.��7oqu���r1��x�����EL���U�\{[U���:P8N�F�n��\b�žh�$�+�rO��˿��<�)����n¦P�~R�Oy^n���3d�BJ�1� [�o�=~���U�n�ceO���ԕUKҪ�Q��=�!��$��/�\(���,��̸rw	�U�M��C��2G?���@���1��3f2�9~vT�1(|��A6*z ���(rx��[���O̇8��Z�M����	�/����b3ݎ��LX�&��ψ%9A���
o��[k�T�Sy/%νȴ���;�uQS*n�Ա^�S��7bmQ8�\��{��Iv�-���}�A)�yq��܊�r��yb�i>�g [��\ f�0Ű��KA��6���4)�54]�њ��vַ�)�j�	+�|U� 
]6:�h�z�/�c7��� �/��w����2������D��֮�˽	'] f�I��A�\q�[�\��CJŻ�۟K;:���=��%��64�S1�Fc�(̯w����������H�3�p�I*-�z���Hd������7(���|c�����Z�D�U�55|��5ZI���K���K���XT�:�������
}�ב��ug�|\��f��AVx�ؗ|��;�ދ#cps&o���plk�+�_�����7��"�"Y�%�/��K��3`���A���>P/�B����gA���M`���Wʳx�D��k.#!N��V��4
i� �H����)��Ha7��N����������m�CQ��?v�bV:��g�m���k�O�\c�쥲%�lq���q�`���gC ���'��G���|8�lo����9�8c;#v�[�K���O�^NBƄz�+q+��o��$��t� ]g0�鉺�{��{��P�aAc���ީ���K�*�d_C�L?�^?^��~$�C.�ЕJV�E�@�)ͱ�y�
��0֟�4�U�����tC!���`;"tP�X }�@z����b˾8pGZ)V�����,q���e[u�b��@�Y�n�r������_� d�/8A=V�g���qUl���_���.X�[Ҁk����n�#sSN$u�n���`!���.�?CtmƠcg��cA�8�T��(e��؅$Z��{�h�3hBh	��x�+�j����e�.@I�p�`-�O,P���]U�ޅ�Ƃ�оq�>wo�.�鲄�8��7Td���FNjo���$oL�.����W�\��v�Rq��ι�ҩ4��G{h�Sꝲ��
"V�#g�66c�"��3O��4wH���g��@$�qE�n�t�	�O*8}�XCͮأ�q�ш�ɇ���SG�+Θ��u�qLGm�B���L'򂟋�a���\2�?S2�Qb�_=�?��