
module nios (
	clk_clk);	

	input		clk_clk;
endmodule
