
module DE0_NANO_SOPC (
	clk_clk);	

	input		clk_clk;
endmodule
