
module CPU (
	clk_clk);	

	input		clk_clk;
endmodule
